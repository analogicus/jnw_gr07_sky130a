*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/temp_to_current_tb_lpe.spi
#else
.include ../../../work/xsch/temp_to_current_tb.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD VDD 0 dc {AVDD}


*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
*.TEMP -40 -20 0 20 40 60 80 100 120

.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 10u 0

dc temp -40 120 20 ; sweep dc operating points vs temp

* tran 1n 10n 1p
write
quit


.endc

.end
