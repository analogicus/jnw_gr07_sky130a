magic
tech sky130A
magscale 1 2
timestamp 1744468687
<< locali >>
rect 5702 8096 9798 8100
rect 5702 7704 9832 8096
rect 8488 7328 8680 7704
rect 9640 7376 9832 7704
rect 8488 4576 8680 6896
rect 9640 4576 9832 6996
rect 8488 3896 8680 4096
rect 9640 3896 9832 4096
rect 8488 3704 9832 3896
rect 4400 -2700 8000 -2000
rect 8480 -2700 8536 -2616
rect 4400 -2900 9500 -2700
rect 4400 -3500 5200 -2900
rect 0 -3739 5200 -3500
rect 6100 -3739 6800 -2900
rect 7700 -3664 8400 -2900
rect 7700 -3739 8461 -3664
rect 0 -3800 5261 -3739
rect 5964 -3800 8536 -3739
rect 9300 -3800 9500 -2900
rect 0 -3900 9500 -3800
rect 0 -7100 100 -3900
rect 4400 -4500 9500 -3900
rect 4400 -5400 5261 -4500
rect 6100 -5339 6800 -4500
rect 6079 -5400 6936 -5339
rect 7700 -5400 8461 -4500
rect 9300 -5400 9500 -4500
rect 4400 -6100 9500 -5400
rect 4400 -6136 5261 -6100
rect 6064 -6121 8461 -6100
rect 4400 -7000 5200 -6136
rect 6100 -7000 6800 -6121
rect 7700 -6136 8461 -6121
rect 7700 -7000 8400 -6136
rect 9300 -7000 9500 -6100
rect 4400 -7075 9500 -7000
rect 4251 -7100 9500 -7075
rect 0 -7400 9500 -7100
rect 0 -7500 5100 -7400
rect 0 -10800 100 -7500
rect 4400 -10800 4900 -7500
<< viali >>
rect 8480 -2616 8536 -2572
rect 364 -4280 604 -4040
rect 3880 -4280 4108 -4040
rect 380 -7880 620 -7640
rect 3868 -7880 4108 -7640
rect 5164 -7880 5404 -7640
rect 8668 -7880 8908 -7640
<< metal1 >>
rect 2304 7904 4296 8096
rect 7072 7904 9064 8096
rect 7072 7404 7264 7904
rect 8744 3532 8808 6932
rect 8872 4304 9064 7904
rect 9256 6404 9448 6996
rect 9256 5296 9448 5596
rect 9256 5098 9448 5104
rect 9256 3896 9448 4296
rect 9256 3698 9448 3704
rect 8168 3468 8808 3532
rect 8168 432 8232 3468
rect 7468 368 8232 432
rect 8168 -968 8232 368
rect 8168 -1032 8568 -968
rect 8632 -1032 8638 -968
rect 4580 -2420 5380 -2180
rect 5620 -2420 5626 -2180
rect 180 -4040 620 -4020
rect 180 -4280 364 -4040
rect 604 -4280 620 -4040
rect 180 -4300 620 -4280
rect 3874 -4040 4114 -4028
rect 4580 -4040 4820 -2420
rect 8468 -2572 8672 -2566
rect 8468 -2616 8480 -2572
rect 8536 -2616 8672 -2572
rect 8468 -2622 8672 -2616
rect 8728 -2622 8734 -2566
rect 5800 -3180 8600 -3100
rect 5580 -3400 8908 -3180
rect 3874 -4280 3880 -4040
rect 4108 -4280 4820 -4040
rect 5400 -3600 9100 -3400
rect 3874 -4292 4114 -4280
rect 180 -7620 420 -4300
rect 5400 -6300 5900 -3600
rect 7180 -4080 7420 -4074
rect 7180 -5020 7420 -4320
rect 8600 -6300 9100 -3600
rect 5400 -6400 9100 -6300
rect 5400 -6500 8908 -6400
rect 5580 -6620 8908 -6500
rect 5900 -6800 8908 -6620
rect 8668 -7620 8908 -6800
rect 180 -7640 640 -7620
rect 180 -7880 380 -7640
rect 620 -7880 640 -7640
rect 180 -7900 640 -7880
rect 3860 -7640 4120 -7620
rect 5140 -7640 5420 -7620
rect 3860 -7880 3868 -7640
rect 4108 -7880 5164 -7640
rect 5404 -7880 5420 -7640
rect 3860 -7900 4120 -7880
rect 5140 -7900 5420 -7880
rect 8660 -7640 8920 -7620
rect 8660 -7880 8668 -7640
rect 8908 -7880 8920 -7640
rect 8660 -7900 8920 -7880
<< via1 >>
rect 9256 5104 9448 5296
rect 9256 3704 9448 3896
rect 8568 -1032 8632 -968
rect 5380 -2420 5620 -2180
rect 8672 -2622 8728 -2566
rect 7180 -4320 7420 -4080
<< metal2 >>
rect 8095 5104 8104 5296
rect 8286 5104 9256 5296
rect 9448 5104 9454 5296
rect 8080 3896 9460 3900
rect 8080 3704 9256 3896
rect 9448 3704 9460 3896
rect 8080 3660 9460 3704
rect 5380 -2180 5620 -2174
rect 5620 -2420 6690 -2180
rect 6920 -2420 6929 -2180
rect 5380 -2426 5620 -2420
rect 8080 -4080 8320 3660
rect 8568 -968 8632 -962
rect 8632 -1032 8776 -968
rect 8832 -1032 8841 -968
rect 8568 -1038 8632 -1032
rect 8672 -2566 8728 -2560
rect 8728 -2622 8872 -2566
rect 8928 -2622 8937 -2566
rect 8672 -2628 8728 -2622
rect 7174 -4320 7180 -4080
rect 7420 -4320 8320 -4080
<< via2 >>
rect 8104 5104 8286 5296
rect 6690 -2420 6920 -2180
rect 8776 -1032 8832 -968
rect 8872 -2622 8928 -2566
<< metal3 >>
rect 8080 5296 8320 5320
rect 8080 5104 8104 5296
rect 8286 5104 8320 5296
rect 6685 -2180 6925 -2175
rect 8080 -2180 8320 5104
rect 8771 -968 8837 -963
rect 8771 -1032 8776 -968
rect 8832 -1032 8837 -968
rect 8771 -1037 8837 -1032
rect 8772 -1632 8836 -1037
rect 6685 -2420 6690 -2180
rect 6920 -2420 8320 -2180
rect 6685 -2425 6925 -2420
rect 8867 -2564 8933 -2561
rect 9062 -2564 9068 -2562
rect 8867 -2566 9068 -2564
rect 8867 -2622 8872 -2566
rect 8928 -2622 9068 -2566
rect 8867 -2624 9068 -2622
rect 8867 -2627 8933 -2624
rect 9062 -2626 9068 -2624
rect 9132 -2626 9138 -2562
<< via3 >>
rect 9068 -2626 9132 -2562
<< metal4 >>
rect 9070 -2561 9130 -2370
rect 9067 -2562 9133 -2561
rect 9067 -2626 9068 -2562
rect 9132 -2626 9133 -2562
rect 9067 -2627 9133 -2626
use amplifier_rev2  amplifier_rev2_0 ../JNW_GR07_SKY130A
timestamp 1744468687
transform 1 0 1000 0 1 -200
box -1600 -3400 7200 8300
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1736794646
transform 1 0 8200 0 1 -5600
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1736794646
transform 1 0 5000 0 1 -7200
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1736794646
transform 1 0 5000 0 1 -5600
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1736794646
transform 1 0 6600 0 1 -7200
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1736794646
transform 1 0 8200 0 1 -7200
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1736794646
transform 1 0 5000 0 1 -4000
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1736794646
transform 1 0 6600 0 1 -4000
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1736794646
transform 1 0 6600 0 1 -5600
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1736794646
transform 1 0 8200 0 1 -4000
box 0 0 1340 1340
use JNWTR_CAPX1  x2 ../JNW_TR_SKY130A
timestamp 1744368984
transform 1 0 8400 0 1 -2400
box 0 0 1080 1080
use JNWATR_PCH_4C5F0  x3 ../JNW_ATR_SKY130A
timestamp 1744368984
transform 1 0 8584 0 1 3928
box -184 -128 1336 928
use JNWTR_RPPO16  x4 ../JNW_TR_SKY130A
timestamp 1744468687
transform 1 0 0 0 1 -7200
box 0 0 4472 3440
use JNWATR_PCH_4C5F0  x5
timestamp 1744368984
transform 1 0 8584 0 1 6728
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  x
timestamp 1744368984
transform 1 0 8584 0 1 5328
box -184 -128 1336 928
use JNWTR_RPPO16  x6
timestamp 1744468687
transform -1 0 4472 0 1 -10800
box 0 0 4472 3440
use JNWTR_RPPO16  x7
timestamp 1744468687
transform -1 0 9272 0 1 -10800
box 0 0 4472 3440
<< labels >>
flabel metal1 9256 6404 9448 6596 0 FreeSans 1600 0 0 0 I_OUT
port 1 nsew
flabel locali 4400 -10800 4900 -10300 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
flabel metal1 2304 7904 2496 8096 0 FreeSans 1600 0 0 0 VDD
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 32656 3440
<< end >>
