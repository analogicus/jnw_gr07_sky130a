* TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/temperature_to_current_tord_lpe.spi
#else
.include ../../../work/xsch/temperature_to_current_tord.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

*
* original code stops, self written code begins ...
*

* fix taken from jnw_gr05
.param vdda = 1.8

*
* self written code stops, original code continues...
*

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
*VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}
*IBP 0 IBPS_5U dc 5u
*V0  IBNS_20U 0 dc 1

*
* original code stops, self written code begins ...
*

VDD VDD_1V8 VSS dc 1.8
V_PTAT I_PTAT VSS dc 0.5 

*
* V_PTAT value of 0.5 is some magic number that was given to us by Carsten
*

*
* self written code stops, original code continues...
*

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
.include ../../../../cpdk/ngspice/ideal_circuits.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
*.probe I(xdut.R1)
*.probe alli
*.option savecurrents
*.save all
.save @r.xdut.r1[i]
.save i(v_ptat)
.save v(v_d1)
.save v(v_ref)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0
*tran 1n 10000n 1p
*.dc TEMP -40 125 10

*write

*
* original code stops, self written code begins ...
*

set fend = .raw
foreach vtemp -40, -35, -30, -25, -20, -15, -10, -5, 0, 5, 10, 15, 20, 25, 30, 35, 40, 45, 50, 55, 60, 65, 70, 75, 80, 85, 90, 95, 100, 105, 110, 115, 120
	option temp=$vtemp
	tran 1n 10u 10n
	write {cicname}_$vtemp$fend
end

*
* self written code stops, original code continues...
*

quit

.endc

.end
