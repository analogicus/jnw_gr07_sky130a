*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/amplifier_lpe.spi
#else
.include ../../../work/xsch/amplifier.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
V0 VDD VSS dc 3.3
V1 Vin+ VSS dc 1 ac 10m 0
*V1 Vin+ VSS sin(1 10mV 1k)
V2 Vin- VSS dc 1

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all
.save v(vin+)
.save v(vout)


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

* optran 0 0 0 1n 1u 0

tran 1n 2m 1p;
* AC analysis from 1Hz to 1GHz with 10 points per decade
* ac dec 10 1k 1Meg
* tran 1n 10n 1p
ac lin 1 1k 1k
write
quit


.endc

.end
