*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/temp_to_current_lpe.spi
#else
.include ../../../work/xsch/temp_to_current.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD  VSS dc {AVDD}
Vmeasure I_OUT point dc 0
Rout point VSS 1k

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all
*.save i(vmeasure)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

*optran 0 0 0 1n 1u 0

*dc temp -40 120 20 ; sweep dc operating points vs temp
*write

set fend = .raw
foreach vtemp -40 -20 0 20 40 60 80 100 120
     option  temp=$vtemp
     tran 10n 5u
     write {cicname}_$vtemp$fend
end

quit


.endc

.end
