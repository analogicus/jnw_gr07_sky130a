magic
tech sky130A
magscale 1 2
timestamp 1744366208
<< locali >>
rect 10044 21096 10336 21176
rect 9988 21090 11332 21096
rect 8562 21044 9132 21054
rect 7788 20852 8556 21044
rect 8736 20862 9132 21044
rect 7788 20676 7980 20852
rect 8940 20672 9132 20862
rect 9988 20910 10110 21090
rect 10290 20910 11332 21090
rect 9988 20904 11332 20910
rect 9988 20884 10336 20904
rect 9988 20676 10180 20884
rect 11140 20676 11332 20904
rect 9988 19376 10180 20196
rect 11140 19328 11332 20196
rect 5918 18100 7264 18340
rect 7492 18100 7496 18340
rect 5906 15032 6740 15120
rect 5879 14976 6740 15032
rect 5906 14880 6740 14976
rect 12800 11880 13620 12120
rect 12800 7180 13620 7420
rect 12800 2880 13620 3120
rect 14183 1683 14218 1914
rect 15585 1683 15620 1914
rect 16985 1683 17020 1914
rect 18385 1683 18420 1914
rect 12800 480 19120 720
rect 14184 283 14219 480
rect 15584 283 15619 480
rect 16984 283 17019 480
rect 18385 283 18420 480
<< viali >>
rect 8556 20852 8736 21044
rect 10110 20910 10290 21090
rect 7264 18100 7492 18340
rect 13874 15374 13926 15426
rect 13780 11764 14020 11992
rect 13786 10686 14014 10914
rect 13780 7180 14020 7408
rect 13786 6086 14014 6314
rect 13780 2580 14020 2808
<< metal1 >>
rect 6924 21204 10296 21396
rect 6267 14854 6334 14860
rect 5667 14787 6267 14854
rect 6267 14781 6334 14787
rect 6924 12304 7116 21204
rect 8556 21056 8748 21204
rect 10104 21176 10296 21204
rect 8550 21044 8748 21056
rect 8550 20852 8556 21044
rect 8736 20852 8748 21044
rect 10044 21096 10336 21176
rect 10044 21090 10596 21096
rect 10044 20910 10110 21090
rect 10290 20910 10596 21090
rect 10044 20904 10596 20910
rect 10044 20884 10336 20904
rect 8550 20840 8748 20852
rect 8556 20524 8748 20840
rect 10372 20504 10564 20904
rect 10756 20596 10948 21296
rect 8172 19896 8364 20260
rect 7604 19753 8364 19896
rect 8812 19832 8876 20132
rect 9104 19832 9288 19836
rect 8812 19768 9288 19832
rect 7587 19704 8364 19753
rect 7258 18652 7498 18658
rect 7258 18340 7498 18412
rect 7258 18100 7264 18340
rect 7492 18100 7498 18340
rect 7258 18088 7498 18100
rect 7587 14854 7654 19704
rect 9104 18796 9288 19768
rect 10244 18796 10308 20152
rect 10372 19104 10564 20396
rect 9096 18604 9102 18796
rect 9294 18608 10308 18796
rect 10868 18768 11632 18832
rect 9294 18604 10296 18608
rect 9524 18504 9716 18604
rect 7261 14787 7267 14854
rect 7334 14787 7837 14854
rect 11568 14852 11632 18768
rect 13268 15426 13938 15432
rect 13268 15374 13874 15426
rect 13926 15374 13938 15426
rect 13268 15368 13938 15374
rect 13268 14852 13332 15368
rect 11568 14788 13332 14852
rect 13768 11992 14032 11998
rect 13768 11764 13780 11992
rect 14020 11764 14032 11992
rect 13768 11758 14032 11764
rect 13780 10914 14020 11758
rect 13780 10686 13786 10914
rect 14014 10686 14020 10914
rect 13780 10674 14020 10686
rect 13768 7408 14032 7414
rect 13768 7180 13780 7408
rect 14020 7180 14032 7408
rect 13768 7174 14032 7180
rect 13780 6314 14020 7174
rect 13780 6086 13786 6314
rect 14014 6086 14020 6314
rect 13780 6074 14020 6086
rect 13768 2808 14032 2814
rect 13768 2580 13780 2808
rect 14020 2580 14032 2808
rect 13768 2574 14032 2580
rect 13780 1620 14020 2574
rect 13780 1380 18720 1620
rect 13780 -280 14020 1380
rect 13780 -520 18720 -280
<< via1 >>
rect 6267 14787 6334 14854
rect 7258 18412 7498 18652
rect 9102 18604 9294 18796
rect 7267 14787 7334 14854
<< metal2 >>
rect 7258 18996 7498 19005
rect 7258 18652 7498 18766
rect 9102 18796 9294 18802
rect 7252 18412 7258 18652
rect 7498 18412 7504 18652
rect 9102 18580 9294 18604
rect 9102 18389 9294 18398
rect 7267 14854 7334 14860
rect 6261 14787 6267 14854
rect 6334 14787 7267 14854
rect 7267 14781 7334 14787
<< via2 >>
rect 7258 18766 7498 18996
rect 9102 18398 9294 18580
<< metal3 >>
rect 7258 19354 7498 19360
rect 7258 19001 7498 19116
rect 7253 18996 7503 19001
rect 7253 18766 7258 18996
rect 7498 18766 7503 18996
rect 7253 18761 7503 18766
rect 8438 18585 8630 19116
rect 8438 18580 9299 18585
rect 8438 18398 9102 18580
rect 9294 18398 9299 18580
rect 8438 18393 9299 18398
<< via3 >>
rect 7258 19116 7498 19354
<< metal4 >>
rect 7257 19354 8532 19355
rect 7257 19116 7258 19354
rect 7498 19116 8532 19354
rect 7257 19115 8532 19116
use amplifier  amplifier_0
timestamp 1744276743
transform 0 -1 15920 1 0 1620
box -3420 2880 17196 9420
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 10084 0 1 18628
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_1
timestamp 1734044400
transform 1 0 10084 0 1 20028
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_2
timestamp 1734044400
transform -1 0 9036 0 -1 20828
box -184 -128 1336 928
use JNWTR_RPPO16  JNWTR_RPPO16_0 ../JNW_TR_SKY130A
timestamp 1744276743
transform 0 -1 16940 1 0 2200
box 0 0 4472 3440
use JNWTR_RPPO16  JNWTR_RPPO16_1
timestamp 1744276743
transform 0 -1 16940 1 0 11400
box 0 0 4472 3440
use JNWTR_RPPO16  JNWTR_RPPO16_2
timestamp 1744276743
transform 0 -1 16940 1 0 6800
box 0 0 4472 3440
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1736794646
transform 1 0 14900 0 1 -800
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1736794646
transform 1 0 13500 0 1 -800
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1736794646
transform 1 0 16300 0 1 -800
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1736794646
transform 1 0 17700 0 1 -800
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1736794646
transform 1 0 13500 0 1 600
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1736794646
transform 1 0 14900 0 1 600
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1736794646
transform 1 0 16300 0 1 600
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1736794646
transform 1 0 17700 0 1 600
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1736794646
transform 1 0 4800 0 1 14100
box 0 0 1340 1340
use JNWTR_CAPX1  x2 ../JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 7880 0 1 18504
box 0 0 1080 1080
<< labels >>
flabel metal1 6924 21204 10296 21396 0 FreeSans 1600 0 0 0 VDD
port 2 nsew
flabel locali 5918 18100 6158 18340 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal1 10756 21104 10948 21296 0 FreeSans 1600 0 0 0 I_OUT
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 32656 3440
<< end >>
