magic
tech sky130A
magscale 1 2
timestamp 1744368116
<< locali >>
rect 22750 23070 22810 23170
rect 12780 22800 13020 22820
rect 12780 22794 14812 22800
rect 12780 22630 14642 22794
rect 14806 22630 14812 22794
rect 12780 22624 14812 22630
rect 19238 22636 19530 22696
rect 12780 18100 13020 22624
rect 19238 21654 19298 22636
rect 21950 21770 22082 21830
rect 19239 20869 19297 21654
rect 19227 20863 19309 20869
rect 19227 20817 19239 20863
rect 19297 20817 19309 20863
rect 19227 20811 19309 20817
rect 22742 20764 22802 20916
rect 18076 20412 18896 20604
rect 19376 20412 20196 20604
rect 20016 20190 20184 20412
rect 20016 20034 20022 20190
rect 20178 20034 20184 20190
rect 20016 19580 20184 20034
rect 22218 19670 22634 19730
rect 18076 19388 18796 19580
rect 19376 19388 20184 19580
rect 20016 18116 20184 19388
rect 22814 19106 23366 19166
rect 21454 18728 22564 18808
rect 21454 18218 21534 18728
rect 26300 16280 27320 16520
rect 19646 15500 20240 15740
rect 26300 13480 26920 13720
rect 26300 11480 26920 11720
rect 18880 480 20220 720
<< viali >>
rect 22750 23170 22810 23230
rect 14642 22630 14806 22794
rect 22082 21770 22130 21830
rect 22742 20916 22802 20964
rect 19239 20817 19297 20863
rect 20022 20034 20178 20190
rect 22170 19670 22218 19730
rect 23366 19106 23426 19166
rect 19418 15500 19646 15740
rect 27172 15472 27227 15527
rect 27172 14173 27227 14228
rect 27086 13186 27314 13414
rect 27080 11888 27320 12116
rect 27080 10980 27320 11208
rect 27086 9686 27314 9914
rect 27080 8764 27320 9004
<< metal1 >>
rect 19070 23291 19130 23330
rect 19070 23230 20250 23291
rect 22750 23250 22810 23730
rect 15914 22800 16090 22806
rect 14630 22794 15914 22800
rect 14630 22630 14642 22794
rect 14806 22630 15914 22794
rect 14630 22624 15914 22630
rect 15914 22618 16090 22624
rect 19070 22436 19130 23230
rect 20230 23170 20250 23230
rect 22730 23230 22830 23250
rect 22730 23170 22750 23230
rect 22810 23170 22830 23230
rect 22730 23150 22830 23170
rect 19064 22430 19136 22436
rect 19064 22370 19070 22430
rect 19130 22370 19136 22430
rect 19064 22364 19136 22370
rect 22076 21830 22136 21842
rect 9906 21612 9912 21788
rect 10088 21612 10094 21788
rect 22076 21770 22082 21830
rect 22130 21770 22170 21830
rect 22230 21770 22236 21830
rect 22076 21758 22136 21770
rect 9912 21212 10088 21612
rect 10750 21328 10756 21520
rect 10948 21328 10954 21520
rect 10756 21104 10948 21328
rect 22730 20964 23024 20970
rect 22730 20916 22742 20964
rect 22802 20916 23024 20964
rect 22730 20910 23024 20916
rect 23084 20910 23090 20970
rect 19227 20863 19309 20869
rect 19227 20817 19239 20863
rect 19297 20817 19309 20863
rect 19227 20811 19309 20817
rect 18068 20284 18932 20348
rect 19239 20291 19297 20811
rect 22164 20730 22224 20736
rect 18016 20028 18936 20196
rect 19320 20190 20190 20196
rect 19320 20034 20022 20190
rect 20178 20034 20190 20190
rect 19320 20028 20190 20034
rect 16195 19964 16407 19974
rect 16195 19772 16204 19964
rect 16396 19772 17696 19964
rect 17996 19772 18896 19964
rect 16195 19762 16407 19772
rect 22164 19730 22224 20670
rect 24554 20040 24560 20280
rect 24800 20040 30580 20280
rect 22164 19670 22170 19730
rect 22218 19670 22224 19730
rect 22164 19658 22224 19670
rect 23324 19166 23516 19236
rect 23324 19106 23366 19166
rect 23426 19106 23516 19166
rect 23324 18418 23516 19106
rect 19412 15740 19652 15752
rect 18862 15500 18868 15740
rect 19108 15500 19418 15740
rect 19646 15500 19652 15740
rect 19412 15488 19652 15500
rect 27166 15527 27233 15539
rect 27166 15472 27172 15527
rect 27227 15472 27233 15527
rect 27166 14854 27233 15472
rect 19600 14788 19606 14852
rect 19670 14788 21614 14852
rect 25267 14787 27233 14854
rect 27166 14228 27233 14787
rect 27166 14173 27172 14228
rect 27227 14173 27233 14228
rect 27166 14161 27233 14173
rect 27080 13414 27320 13426
rect 27080 13186 27086 13414
rect 27314 13186 27320 13414
rect 27080 12122 27320 13186
rect 27068 12116 27332 12122
rect 27068 11888 27080 12116
rect 27320 11888 27332 12116
rect 27068 11882 27332 11888
rect 27068 11208 27332 11214
rect 27068 10980 27080 11208
rect 27320 10980 27332 11208
rect 27068 10974 27332 10980
rect 27080 9914 27320 10974
rect 27080 9686 27086 9914
rect 27314 9686 27320 9914
rect 27080 9674 27320 9686
rect 27070 9004 27340 9030
rect 25980 8764 27080 9004
rect 27320 8764 27340 9004
rect 26700 8320 26940 8764
rect 27070 8750 27340 8764
rect 30340 8320 30580 20040
rect 26700 8080 30580 8320
<< via1 >>
rect 15914 22624 16090 22800
rect 19070 22370 19130 22430
rect 9912 21612 10088 21788
rect 22170 21770 22230 21830
rect 10756 21328 10948 21520
rect 23024 20910 23084 20970
rect 22164 20670 22224 20730
rect 16204 19772 16396 19964
rect 24560 20040 24800 20280
rect 18868 15500 19108 15740
rect 19606 14788 19670 14852
<< metal2 >>
rect 16999 22800 17165 22804
rect 15908 22624 15914 22800
rect 16090 22795 17170 22800
rect 16090 22629 16999 22795
rect 17165 22629 17170 22795
rect 16090 22624 17170 22629
rect 16999 22620 17165 22624
rect 18855 22430 18935 22435
rect 19064 22430 19136 22436
rect 18855 22370 18870 22430
rect 18926 22370 19070 22430
rect 19130 22370 19136 22430
rect 18855 22365 18935 22370
rect 19064 22364 19136 22370
rect 9917 22260 10083 22264
rect 9912 22255 10088 22260
rect 9912 22089 9917 22255
rect 10083 22089 10088 22255
rect 9912 21788 10088 22089
rect 9912 21606 10088 21612
rect 22170 21830 22230 21836
rect 10756 21520 10948 21526
rect 10948 21510 12236 21520
rect 10948 21328 12222 21510
rect 12418 21328 12427 21520
rect 10756 21322 10948 21328
rect 12222 21319 12414 21328
rect 22170 21030 22230 21770
rect 22164 20970 22230 21030
rect 23024 20970 23084 20976
rect 22164 20730 22224 20970
rect 23084 20910 23198 20970
rect 23254 20910 23263 20970
rect 23024 20904 23084 20910
rect 22158 20670 22164 20730
rect 22224 20670 22230 20730
rect 23338 20268 23562 20282
rect 24560 20280 24800 20286
rect 23332 20263 24560 20268
rect 23332 20097 23377 20263
rect 23543 20097 24560 20263
rect 23332 20092 24560 20097
rect 23332 20078 23562 20092
rect 24560 20034 24800 20040
rect 16195 19964 16407 19974
rect 16195 19772 16204 19964
rect 16396 19772 16407 19964
rect 16195 19762 16407 19772
rect 16204 19491 16396 19762
rect 16191 19486 16401 19491
rect 16191 19304 16204 19486
rect 16396 19304 16401 19486
rect 16191 19295 16401 19304
rect 16191 19292 16400 19295
rect 18868 16164 19108 16173
rect 18868 15740 19108 15934
rect 18868 15494 19108 15500
rect 19606 14852 19670 14858
rect 17777 14788 17786 14852
rect 17842 14788 19606 14852
rect 19606 14782 19670 14788
<< via2 >>
rect 16999 22629 17165 22795
rect 18870 22370 18926 22430
rect 9917 22089 10083 22255
rect 12236 21510 12418 21520
rect 12222 21328 12418 21510
rect 23198 20910 23254 20970
rect 23377 20097 23543 20263
rect 16204 19304 16396 19486
rect 18868 15934 19108 16164
rect 17786 14788 17842 14852
<< metal3 >>
rect 16994 22795 19788 22800
rect 16994 22629 16999 22795
rect 17165 22629 19788 22795
rect 16994 22624 19788 22629
rect 23084 22624 23928 22800
rect 18855 22430 18935 22435
rect 18855 22370 18870 22430
rect 18926 22370 18935 22430
rect 18855 22365 18935 22370
rect 18868 22260 18928 22365
rect 9912 22255 19788 22260
rect 9912 22089 9917 22255
rect 10083 22089 19788 22255
rect 9912 22084 19788 22089
rect 23084 22084 23548 22260
rect 12231 21520 12423 21525
rect 12231 21515 12236 21520
rect 12217 21510 12236 21515
rect 12217 21328 12222 21510
rect 12418 21328 12423 21520
rect 12217 21323 12423 21328
rect 12231 18840 12423 21323
rect 23193 20970 23259 20975
rect 23372 20970 23548 22084
rect 23193 20910 23198 20970
rect 23254 20910 23548 20970
rect 23193 20905 23259 20910
rect 23372 20263 23548 20910
rect 23372 20100 23377 20263
rect 22828 20097 23377 20100
rect 23543 20097 23548 20263
rect 22828 19924 23548 20097
rect 23752 19560 23928 22624
rect 16184 19486 16401 19491
rect 16184 19304 16204 19486
rect 16396 19304 16401 19486
rect 22828 19384 23928 19560
rect 16184 19295 16401 19304
rect 16184 19292 16400 19295
rect 16204 18840 16396 19292
rect 12231 18648 16396 18840
rect 16204 17344 16396 18648
rect 16204 17152 17916 17344
rect 17782 14857 17846 17152
rect 18863 16164 19412 16169
rect 18863 15934 18868 16164
rect 19108 15934 19412 16164
rect 18863 15929 19412 15934
rect 19650 15929 19656 16169
rect 17781 14852 17847 14857
rect 17781 14788 17786 14852
rect 17842 14788 17847 14852
rect 17781 14783 17847 14788
<< via3 >>
rect 19412 15929 19650 16169
<< metal4 >>
rect 19411 16169 19651 16966
rect 19411 15929 19412 16169
rect 19650 15929 19651 16169
rect 19411 15928 19651 15929
use amplifier  amplifier_1
timestamp 1744276743
transform 0 1 17120 1 0 1620
box -3420 2880 17196 9420
use JNWATR_NCH_2C1F2  JNWATR_NCH_2C1F2_1 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 0 1 17428 -1 0 20508
box -184 -128 1208 928
use JNWATR_NCH_2C1F2  JNWATR_NCH_2C1F2_2
timestamp 1734044400
transform 0 1 18728 -1 0 20508
box -184 -128 1208 928
use JNWTR_BFX1_CV  JNWTR_BFX1_CV_1 ../JNW_TR_SKY130A
timestamp 1744366080
transform 0 -1 23004 1 0 18754
box -150 -120 2130 600
use JNWTR_DFRNQNX1_CV  JNWTR_DFRNQNX1_CV_1 ../JNW_TR_SKY130A
timestamp 1744366080
transform 0 -1 23260 -1 0 23430
box -150 -120 2130 3960
use JNWTR_RPPO4  JNWTR_RPPO4_1 ../JNW_TR_SKY130A
timestamp 1744276743
transform 0 -1 30240 -1 0 14680
box 0 0 1880 3440
use JNWTR_RPPO4  JNWTR_RPPO4_2
timestamp 1744276743
transform 0 -1 30240 -1 0 12480
box 0 0 1880 3440
use JNWTR_RPPO4  JNWTR_RPPO4_3
timestamp 1744276743
transform 0 -1 30240 -1 0 10280
box 0 0 1880 3440
use JNWTR_RPPO4  JNWTR_RPPO4_4
timestamp 1744276743
transform 0 -1 30240 -1 0 16880
box 0 0 1880 3440
use temp_to_current  temp_to_current_1
timestamp 1744366208
transform 1 0 0 0 1 0
box 4800 -1800 19120 21396
<< labels >>
flabel metal3 12412 22084 12588 22260 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel metal1 22750 23670 22810 23730 0 FreeSans 1600 0 0 0 CLK
port 3 nsew
flabel locali 13672 22624 13848 22800 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel locali 19239 20863 19297 22696 0 FreeSans 1600 0 0 0 PWM
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 62144 3840
<< end >>
