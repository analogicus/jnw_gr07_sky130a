magic
tech sky130A
magscale 1 2
timestamp 1744010837
<< error_s >>
rect 4700 7700 6220 7710
rect 6500 7700 8020 7710
rect 8300 7700 9820 7710
rect 13300 6600 13310 8120
rect 16492 6688 16498 6700
rect 16702 6688 16708 6700
rect 16504 6676 16516 6682
rect 16684 6676 16696 6682
rect 4700 6400 6220 6410
rect 6500 6400 8020 6410
rect 8300 6400 9820 6410
rect 4700 5100 6220 5110
rect 6500 5100 8020 5110
rect 8300 5100 9820 5110
rect 13300 4500 13310 6020
rect 15362 5612 15368 5618
rect 15432 5612 15438 5618
rect 15368 5606 15374 5612
rect 15426 5606 15432 5612
rect 3862 4146 3910 4152
rect 4090 4146 4102 4152
rect 4114 4146 4130 4174
rect 3862 4140 3878 4146
rect 4074 4112 4096 4146
rect 4102 4140 4130 4146
<< locali >>
rect -2780 9380 16720 9420
rect -3420 9180 16720 9380
rect -3420 3120 -3180 9180
rect 16480 8032 16720 9180
rect 4788 7204 4980 7980
rect 4789 5905 4979 7204
rect 5940 7176 6132 7996
rect 6588 7176 6780 7996
rect 7740 7176 7932 7996
rect 8388 7176 8580 7996
rect 9540 7104 9732 7980
rect 11984 7840 12296 8032
rect 12804 7840 13596 8032
rect 15176 7840 15696 8032
rect 16176 7840 16516 8032
rect 16696 7880 16720 8032
rect 10288 6804 10300 6996
rect 5940 5876 6132 6696
rect 6588 5876 6780 6696
rect 7740 5876 7932 6696
rect 8388 5876 8580 6696
rect 9540 5876 9732 6696
rect 10288 6576 10480 6804
rect 11440 6576 11632 6816
rect 11984 6688 12296 6880
rect 12776 6688 13596 6880
rect 15176 6688 15696 6880
rect 16176 6688 16504 6880
rect 11984 5740 12296 5932
rect 12776 5740 13596 5932
rect 15176 5740 15696 5932
rect 16128 5740 16516 5932
rect 4788 4504 4980 5380
rect 5940 4528 6132 5496
rect 6588 4576 6780 5396
rect 7740 4576 7932 5396
rect 8388 4576 8580 5396
rect 9540 4576 9732 5396
rect 11984 4588 12280 4780
rect 12776 4588 13596 4780
rect 15176 4588 15696 4780
rect 16176 4588 16516 4780
rect 16696 4588 16720 4720
rect 192 3120 432 4356
rect 4788 3796 4980 4080
rect 5940 3796 6132 4080
rect 6588 3796 6780 4080
rect 7740 3796 7932 4080
rect 8388 3796 8580 4080
rect 9540 3796 9732 4080
rect 16480 3120 16720 4588
rect -3420 2880 16720 3120
<< viali >>
rect 4788 8488 4980 8668
rect 5940 8488 6132 8668
rect 6588 8488 6780 8668
rect 7740 8488 7932 8668
rect 8388 8488 8580 8668
rect 9540 8488 9732 8668
rect 192 7632 432 7860
rect 3862 7662 4102 7890
rect 11804 7840 11984 8032
rect 16516 7840 16696 8032
rect 10300 6804 10480 6996
rect 11440 6816 11632 6996
rect 11804 6688 11984 6880
rect 16504 6688 16696 6880
rect 11804 5740 11984 5932
rect 16516 5740 16696 5932
rect 11804 4588 11984 4780
rect 16516 4588 16696 4780
rect 3862 4146 4102 4374
<< metal1 >>
rect 4788 8804 10896 8996
rect 4788 8674 4980 8804
rect 4776 8668 4992 8674
rect 180 8280 4102 8520
rect 4776 8488 4788 8668
rect 4980 8488 4992 8668
rect 4776 8482 4992 8488
rect 5268 8532 5332 8538
rect 5268 8462 5332 8468
rect 5556 8324 5748 8804
rect 5940 8674 6132 8804
rect 6588 8674 6780 8804
rect 5928 8668 6144 8674
rect 5812 8532 5876 8612
rect 5806 8468 5812 8532
rect 5876 8468 5882 8532
rect 5928 8488 5940 8668
rect 6132 8488 6144 8668
rect 5928 8482 6144 8488
rect 6576 8668 6792 8674
rect 6576 8488 6588 8668
rect 6780 8488 6792 8668
rect 6576 8482 6792 8488
rect 7068 8532 7132 8538
rect 5812 8368 5876 8468
rect 7068 8462 7132 8468
rect 7356 8304 7548 8804
rect 7740 8674 7932 8804
rect 8388 8674 8580 8804
rect 7728 8668 7944 8674
rect 7606 8468 7612 8532
rect 7676 8468 7682 8532
rect 7728 8488 7740 8668
rect 7932 8488 7944 8668
rect 7728 8482 7944 8488
rect 8376 8668 8592 8674
rect 8376 8488 8388 8668
rect 8580 8488 8592 8668
rect 8376 8482 8592 8488
rect 8868 8532 8932 8538
rect 7612 8368 7676 8468
rect 8868 8462 8932 8468
rect 9156 8324 9348 8804
rect 9540 8674 9732 8804
rect 9528 8668 9744 8674
rect 9406 8468 9412 8532
rect 9476 8468 9482 8532
rect 9528 8488 9540 8668
rect 9732 8488 9744 8668
rect 9528 8482 9744 8488
rect 9412 8368 9476 8468
rect 192 7866 432 8280
rect 3862 7896 4102 8280
rect 3850 7890 4114 7896
rect 180 7860 444 7866
rect 180 7632 192 7860
rect 432 7632 444 7860
rect 3850 7662 3862 7890
rect 4102 7662 4114 7890
rect 3850 7656 4114 7662
rect 180 7626 444 7632
rect 5172 7232 5364 7996
rect 5172 7168 5268 7232
rect 5332 7168 5364 7232
rect 5172 7096 5364 7168
rect 5556 7024 5748 8096
rect 5812 7232 5876 7932
rect 6972 7232 7164 8060
rect 5806 7168 5812 7232
rect 5876 7168 5882 7232
rect 6972 7168 7068 7232
rect 7132 7168 7164 7232
rect 6972 7104 7164 7168
rect 7356 7004 7548 8132
rect 7612 7232 7676 7932
rect 8772 7232 8964 8060
rect 7606 7168 7612 7232
rect 7676 7168 7682 7232
rect 8772 7168 8868 7232
rect 8932 7168 8964 7232
rect 7612 7068 7676 7168
rect 8772 7104 8964 7168
rect 9156 7104 9348 8132
rect 9412 7232 9476 7932
rect 9406 7168 9412 7232
rect 9476 7168 9482 7232
rect 9412 7068 9476 7168
rect 10294 6996 10486 7008
rect 10672 6996 10864 8804
rect 11798 8032 11990 8044
rect 11798 7840 11804 8032
rect 11984 7840 11990 8032
rect 11798 7648 11990 7840
rect 13167 7776 13234 8333
rect 16510 8032 16702 8044
rect 16510 7996 16516 8032
rect 16504 7840 16516 7996
rect 16696 7840 16702 8032
rect 16504 7828 16702 7840
rect 12824 7712 13532 7776
rect 13167 7711 13234 7712
rect 11798 7456 12432 7648
rect 12604 7456 13732 7648
rect 14304 7456 14760 7648
rect 15004 7456 15796 7648
rect 11798 7404 11996 7456
rect 11428 6996 11644 7002
rect 5172 5932 5364 6796
rect 5172 5868 5268 5932
rect 5332 5868 5364 5932
rect 5172 5796 5364 5868
rect 5556 5724 5748 6796
rect 5812 6332 5876 6612
rect 5806 6268 5812 6332
rect 5876 6268 5882 6332
rect 5812 5932 5876 6268
rect 6972 5932 7164 6760
rect 5806 5868 5812 5932
rect 5876 5868 5882 5932
rect 6972 5868 7068 5932
rect 7132 5868 7164 5932
rect 5812 5768 5876 5868
rect 6972 5804 7164 5868
rect 7356 5704 7548 6832
rect 10294 6804 10300 6996
rect 10480 6816 11440 6996
rect 11632 6816 11644 6996
rect 11804 6892 11996 7404
rect 14304 7264 14496 7456
rect 16504 7264 16696 7828
rect 12696 7072 13696 7264
rect 13996 7072 14496 7264
rect 15024 7072 15896 7264
rect 16004 7072 16696 7264
rect 10480 6810 11644 6816
rect 11798 6880 11996 6892
rect 10480 6804 11596 6810
rect 7612 6332 7676 6632
rect 7612 5932 7676 6268
rect 8772 5932 8964 6760
rect 7606 5868 7612 5932
rect 7676 5868 7682 5932
rect 8772 5868 8868 5932
rect 8932 5868 8964 5932
rect 7612 5768 7676 5868
rect 8772 5804 8964 5868
rect 9156 5724 9348 6796
rect 10294 6792 10486 6804
rect 9412 6332 9476 6632
rect 9412 5932 9476 6268
rect 10544 6332 10608 6338
rect 10672 6304 10864 6804
rect 11798 6688 11804 6880
rect 11984 6688 11996 6880
rect 11798 6676 11996 6688
rect 11804 6396 11996 6676
rect 10544 6164 10608 6268
rect 11056 6204 11996 6396
rect 14304 6396 14496 7072
rect 15168 6944 15368 7008
rect 15432 6944 15732 7008
rect 16504 6886 16696 7072
rect 16498 6880 16702 6886
rect 16498 6688 16504 6880
rect 16696 6688 16702 6880
rect 16498 6682 16702 6688
rect 14304 6204 17196 6396
rect 11056 6004 11248 6204
rect 11804 5944 11996 6204
rect 11798 5932 11996 5944
rect 9406 5868 9412 5932
rect 9476 5868 9482 5932
rect 11798 5740 11804 5932
rect 11984 5740 11996 5932
rect 11798 5728 11996 5740
rect 5172 4632 5364 5496
rect 5172 4568 5268 4632
rect 5332 4568 5364 4632
rect 5172 4496 5364 4568
rect 5556 4424 5748 5496
rect 5812 4632 5876 5332
rect 6972 4632 7164 5496
rect 5806 4568 5812 4632
rect 5876 4568 5882 4632
rect 6972 4568 7068 4632
rect 7132 4568 7164 4632
rect 5812 4468 5876 4568
rect 6972 4404 7164 4568
rect 7356 4424 7548 5496
rect 7612 4632 7676 5332
rect 8772 4632 8964 5396
rect 7606 4568 7612 4632
rect 7676 4568 7682 4632
rect 8772 4568 8868 4632
rect 8932 4568 8964 4632
rect 7612 4468 7676 4568
rect 8772 4496 8964 4568
rect 9156 4424 9348 5496
rect 9412 4632 9476 5332
rect 11804 5196 11996 5728
rect 16510 5932 16702 5944
rect 16510 5740 16516 5932
rect 16696 5740 16702 5932
rect 14304 5676 14496 5696
rect 14304 5612 14652 5676
rect 15168 5612 15368 5676
rect 15432 5612 15732 5676
rect 14304 5548 14496 5612
rect 16510 5548 16702 5740
rect 12696 5356 13696 5548
rect 13904 5356 14496 5548
rect 15004 5356 15796 5548
rect 16004 5356 16702 5548
rect 11798 5164 11996 5196
rect 14304 5164 14496 5356
rect 11798 4972 12496 5164
rect 12704 4972 13732 5164
rect 14304 4972 14796 5164
rect 15096 4972 15796 5164
rect 11798 4780 11990 4972
rect 12768 4844 13532 4908
rect 9406 4568 9412 4632
rect 9476 4568 9482 4632
rect 11798 4588 11804 4780
rect 11984 4588 11990 4780
rect 11798 4576 11990 4588
rect 3850 4374 4114 4380
rect 3850 4140 3862 4374
rect 3904 3496 4096 4146
rect 4102 4140 4114 4374
rect 13168 4268 13232 4844
rect 16510 4780 16702 5356
rect 16510 4588 16516 4780
rect 16696 4588 16702 4780
rect 16510 4576 16702 4588
rect 5172 3496 5364 4196
rect 6972 3496 7164 4160
rect 8772 3496 8964 4160
rect 3904 3304 8996 3496
<< via1 >>
rect 5268 8468 5332 8532
rect 5812 8468 5876 8532
rect 7068 8468 7132 8532
rect 7612 8468 7676 8532
rect 8868 8468 8932 8532
rect 9412 8468 9476 8532
rect 5268 7168 5332 7232
rect 5812 7168 5876 7232
rect 7068 7168 7132 7232
rect 7612 7168 7676 7232
rect 8868 7168 8932 7232
rect 9412 7168 9476 7232
rect 5268 5868 5332 5932
rect 5812 6268 5876 6332
rect 5812 5868 5876 5932
rect 7068 5868 7132 5932
rect 7612 6268 7676 6332
rect 7612 5868 7676 5932
rect 8868 5868 8932 5932
rect 9412 6268 9476 6332
rect 10544 6268 10608 6332
rect 15368 6944 15432 7008
rect 9412 5868 9476 5932
rect 5268 4568 5332 4632
rect 5812 4568 5876 4632
rect 7068 4568 7132 4632
rect 7612 4568 7676 4632
rect 8868 4568 8932 4632
rect 15368 5612 15432 5676
rect 9412 4568 9476 4632
<< metal2 >>
rect 5812 8532 5876 8538
rect 7612 8532 7676 8538
rect 9412 8532 9476 8538
rect 5262 8468 5268 8532
rect 5332 8468 5812 8532
rect 7062 8468 7068 8532
rect 7132 8468 7612 8532
rect 8862 8468 8868 8532
rect 8932 8468 9412 8532
rect 5812 8462 5876 8468
rect 7612 8462 7676 8468
rect 9412 8462 9476 8468
rect 5812 7232 5876 7238
rect 7612 7232 7676 7238
rect 9412 7232 9476 7238
rect 5262 7168 5268 7232
rect 5332 7168 5812 7232
rect 7062 7168 7068 7232
rect 7132 7168 7612 7232
rect 8862 7168 8868 7232
rect 8932 7168 9412 7232
rect 5812 7162 5876 7168
rect 7612 7162 7676 7168
rect 9412 7162 9476 7168
rect 15368 7008 15432 7014
rect 5812 6332 5876 6338
rect 5876 6268 7612 6332
rect 7676 6268 9412 6332
rect 9476 6268 10544 6332
rect 10608 6268 10632 6332
rect 5812 6262 5876 6268
rect 5812 5932 5876 5938
rect 7612 5932 7676 5938
rect 9412 5932 9476 5938
rect 5262 5868 5268 5932
rect 5332 5868 5812 5932
rect 7062 5868 7068 5932
rect 7132 5868 7612 5932
rect 8862 5868 8868 5932
rect 8932 5868 9412 5932
rect 5812 5862 5876 5868
rect 7612 5862 7676 5868
rect 9412 5862 9476 5868
rect 15368 5676 15432 6944
rect 5812 4632 5876 4638
rect 7612 4632 7676 4638
rect 9412 4632 9476 4638
rect 5262 4568 5268 4632
rect 5332 4568 5812 4632
rect 7062 4568 7068 4632
rect 7132 4568 7612 4632
rect 8862 4568 8868 4632
rect 8932 4568 9412 4632
rect 5812 4562 5876 4568
rect 7612 4562 7676 4568
rect 9412 4562 9476 4568
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 0 -1 15328 1 0 6784
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1734044400
transform 0 1 15528 -1 0 5836
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2
timestamp 1734044400
transform 0 1 14528 -1 0 5836
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3
timestamp 1734044400
transform 0 -1 16428 1 0 6784
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform -1 0 9636 0 -1 6028
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_1
timestamp 1734044400
transform -1 0 7836 0 -1 8628
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_2
timestamp 1734044400
transform -1 0 7836 0 -1 4728
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_3
timestamp 1734044400
transform -1 0 6036 0 -1 8628
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_4
timestamp 1734044400
transform -1 0 6036 0 -1 6028
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_5
timestamp 1734044400
transform -1 0 6036 0 -1 4728
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_6
timestamp 1734044400
transform -1 0 9636 0 -1 8628
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_7
timestamp 1734044400
transform -1 0 7836 0 -1 7328
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_8
timestamp 1734044400
transform -1 0 7836 0 -1 6028
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_9
timestamp 1734044400
transform -1 0 9636 0 -1 7328
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_10
timestamp 1734044400
transform -1 0 9636 0 -1 4728
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_11
timestamp 1734044400
transform 0 1 12128 -1 0 7936
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_12
timestamp 1734044400
transform 0 -1 14228 1 0 4684
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_13
timestamp 1734044400
transform 0 -1 12928 1 0 4684
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_14
timestamp 1734044400
transform 0 1 13428 -1 0 7936
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_15
timestamp 1734044400
transform -1 0 6036 0 -1 7328
box -184 -128 1336 928
use JNWTR_RPPO16  x1 ../JNW_TR_SKY130A
timestamp 1743348313
transform 0 1 942 -1 0 8254
box 0 0 4472 3440
use JNWTR_RPPO16  x4
timestamp 1743348313
transform 0 1 -2728 1 0 3752
box 0 0 4472 3440
use JNWATR_PCH_4C5F0  x5
timestamp 1734044400
transform 1 0 10384 0 1 5928
box -184 -128 1336 928
<< labels >>
flabel metal1 6204 8804 6396 8996 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel metal1 13168 4268 13232 4332 0 FreeSans 1600 0 0 0 VINP
port 2 nsew
flabel metal1 13167 8266 13234 8333 0 FreeSans 1600 0 0 0 VINN
port 3 nsew
flabel metal1 17004 6204 17196 6396 0 FreeSans 1600 0 0 0 VOUT
port 4 nsew
flabel locali 880 2880 1120 3120 0 FreeSans 1600 0 0 0 VSS
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 14704 3440
<< end >>
