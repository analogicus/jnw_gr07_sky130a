** sch_path: /home/ranerhei/pro/aicex/ip/jnw_gr07_sky130a/design/JNW_GR07_SKY130A/amplifier_tb.sch
**.subckt amplifier_tb
x1 Vdd_tb Vin+_tb Vin-_tb Vout_tb 0 amplifier
V1 Vin+_tb 0 1
V2 Vin-_tb 0 0.9
V3 Vdd_tb 0 3
C1 Vout_tb 0 10p m=1
**** begin user architecture code



.param mc_mm_switch=0
.param mc_pr_switch=0
.include ~/pro/aicex/ip/jnw_sv_sky130a/design/JNW_SV_SKY130A/simulation/tt.spi
* Options:
.option savecurrents
.option gmin=1e-15
.save all
.control
optran 0 0 0 10n 10u 0
op
write amplifier_tb.raw
exit
.endc
.end


**** end user architecture code
**.ends

* expanding   symbol:  JNW_GR07_SKY130A/amplifier.sym # of pins=5
** sym_path: /home/ranerhei/pro/aicex/ip/jnw_gr07_sky130a/design/JNW_GR07_SKY130A/amplifier.sym
** sch_path: /home/ranerhei/pro/aicex/ip/jnw_gr07_sky130a/design/JNW_GR07_SKY130A/amplifier.sch
.subckt amplifier VDD Vin+ Vin- Vout VSS
*.ipin Vin+
*.ipin Vin-
*.ipin VDD
*.ipin VSS
*.opin Vout
x1 net1 net1 VSS VSS JNWATR_NCH_4C5F0
x2 Vout net1 VSS VSS JNWATR_NCH_4C5F0
x3 net1 Vin+ net2 VDD JNWATR_PCH_4C5F0
x4 Vout Vin- net2 VDD JNWATR_PCH_4C5F0
x5 VDD net2 VSS JNWTR_RES2
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym # of pins=4
** sym_path: /home/ranerhei/pro/aicex/ip/jnw_gr07_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym
** sch_path: /home/ranerhei/pro/aicex/ip/jnw_gr07_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sch
.subckt JNWATR_NCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym # of pins=4
** sym_path: /home/ranerhei/pro/aicex/ip/jnw_gr07_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym
** sch_path: /home/ranerhei/pro/aicex/ip/jnw_gr07_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sch
.subckt JNWATR_PCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES2.sym # of pins=3
** sym_path: /home/ranerhei/pro/aicex/ip/jnw_gr07_sky130a/design/JNW_TR_SKY130A/JNWTR_RES2.sym
** sch_path: /home/ranerhei/pro/aicex/ip/jnw_gr07_sky130a/design/JNW_TR_SKY130A/JNWTR_RES2.sch
.subckt JNWTR_RES2 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 P INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends

.end
