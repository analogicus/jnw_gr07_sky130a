magic
tech sky130A
magscale 1 2
timestamp 1744468687
<< locali >>
rect -1500 8290 5200 8300
rect -1500 8110 1310 8290
rect 1490 8110 5200 8290
rect -1500 8096 5200 8110
rect -1512 7904 5232 8096
rect -1512 7528 -1320 7904
rect -360 7528 480 7904
rect 1440 7528 2280 7904
rect 3240 7528 4080 7904
rect 5040 7528 5232 7904
rect -200 7096 400 7528
rect 1600 7096 2200 7528
rect 3400 7096 4000 7528
rect -1512 4704 -1320 7096
rect -360 4704 480 7096
rect 1440 4704 2280 7096
rect 3240 4704 4080 7096
rect 5040 6596 5232 7096
rect 5040 6404 7032 6596
rect 5040 6128 5880 6404
rect 6840 6128 7032 6404
rect 5040 5496 5800 6128
rect 6840 5496 7032 5696
rect 5040 5304 7032 5496
rect 5040 4704 5232 5304
rect -1512 4096 -1320 4296
rect -200 4096 400 4704
rect 1600 4096 2200 4704
rect 3400 4096 4000 4704
rect 5040 4096 5232 4296
rect -1512 3904 5232 4096
rect -1000 300 -900 3600
rect 3888 3304 6316 3496
rect 6496 3304 7032 3496
rect 3888 2928 4080 3304
rect 5040 2928 5880 3304
rect 6840 2928 7032 3304
rect 5200 2496 5800 2928
rect 3888 1504 4080 2496
rect 5040 1528 5880 2496
rect 6840 1528 7032 2496
rect 5040 1504 5800 1528
rect 3888 896 4080 1096
rect 5200 896 5800 1504
rect 6840 896 7032 1096
rect 3888 704 7032 896
rect 3888 400 7032 496
rect 3400 304 7032 400
rect 3400 300 4080 304
rect -1000 0 4080 300
rect -1000 -3300 -900 0
rect 3400 -72 4080 0
rect 5040 -72 5880 304
rect 6840 -72 7032 304
rect 2868 -480 3108 -80
rect 3400 -504 4000 -72
rect 5200 -504 5800 -72
rect 3400 -1096 4080 -504
rect 5040 -1096 5880 -504
rect 6840 -1096 7032 -504
rect 3400 -1504 4000 -1096
rect 3400 -1704 4080 -1504
rect 5200 -1704 5800 -1096
rect 6840 -1704 7032 -1504
rect 3400 -1896 5304 -1704
rect 5484 -1896 7032 -1704
rect 3400 -3300 3900 -1896
rect -1000 -3400 3900 -3300
<< viali >>
rect 1310 8110 1490 8290
rect -636 3120 -396 3360
rect 2868 3120 3108 3360
rect 6316 3304 6496 3496
rect -636 -480 -396 -240
rect 5304 -1896 5484 -1704
<< metal1 >>
rect -1128 8290 6272 8296
rect -1128 8110 1310 8290
rect 1490 8110 6272 8290
rect -1128 8104 6272 8110
rect -1128 7304 -936 8104
rect -1256 4768 -1192 7232
rect -1128 4504 -936 7296
rect -744 4696 -552 7096
rect -1256 3896 -1192 4232
rect -744 3896 -552 4360
rect 544 3896 608 7632
rect 672 7304 864 8104
rect 672 4504 864 7296
rect 1054 4694 1250 7098
rect 1056 3896 1248 4496
rect 2344 3896 2408 7632
rect 2472 7304 2664 8104
rect 2472 4504 2664 7296
rect 2856 4560 3048 7096
rect 2856 3896 3048 4496
rect 4144 3896 4208 7632
rect 4272 7304 4464 8104
rect 4272 4504 4464 7296
rect 4656 4696 4848 7096
rect 4656 3896 4848 4360
rect 5880 3896 6008 6264
rect 6072 5904 6264 8104
rect -1296 3768 6008 3896
rect -1296 3704 5996 3768
rect 2868 3380 3108 3704
rect 6456 3508 6648 5896
rect 6310 3496 6648 3508
rect -920 3360 -380 3380
rect -920 3120 -636 3360
rect -396 3120 -380 3360
rect -920 3100 -380 3120
rect 2840 3360 3140 3380
rect 2840 3120 2868 3360
rect 3108 3120 3140 3360
rect 4272 3304 6316 3496
rect 6496 3304 6656 3496
rect 2840 3100 3140 3120
rect 4144 3232 4208 3238
rect -920 -220 -680 3100
rect 4144 1568 4208 3168
rect 4272 2704 4464 3304
rect 5944 3232 6008 3238
rect 4272 1304 4464 2696
rect 4656 1496 4848 2496
rect 5944 1368 6008 3168
rect 6072 2704 6264 3304
rect 6310 3292 6502 3304
rect 6072 1304 6264 2696
rect 6456 1304 6648 2696
rect 4656 696 4848 1296
rect 4104 504 6096 696
rect 4144 -32 4208 504
rect -920 -240 -380 -220
rect -920 -480 -636 -240
rect -396 -480 -380 -240
rect 4656 -296 4848 504
rect 5944 -32 6008 504
rect 6456 -96 6648 1296
rect -920 -500 -380 -480
rect 4144 -1032 4208 -568
rect 4272 -1296 4464 -304
rect 4656 -1096 4848 -304
rect 5944 -1032 6008 -568
rect 6072 -1176 6264 -304
rect 6456 -1104 6648 -504
rect 4272 -1706 4464 -1304
rect 5298 -1704 5490 -1692
rect 6072 -1704 6264 -1304
rect 5116 -1706 5304 -1704
rect 4272 -1894 5304 -1706
rect 4272 -1896 4464 -1894
rect 5116 -1896 5304 -1894
rect 5484 -1896 6264 -1704
rect 5298 -1908 5490 -1896
<< via1 >>
rect 4144 3168 4208 3232
rect 5944 3168 6008 3232
<< metal2 >>
rect 4144 3632 4208 3641
rect 4144 3232 4208 3576
rect 4138 3168 4144 3232
rect 4208 3168 4214 3232
rect 5938 3168 5944 3232
rect 6008 3168 7200 3232
<< via2 >>
rect 4144 3576 4208 3632
<< metal3 >>
rect 4139 3636 4213 3637
rect 4139 3632 7198 3636
rect 4139 3576 4144 3632
rect 4208 3576 7198 3632
rect 4139 3572 7198 3576
rect 4139 3571 4213 3572
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1744368984
transform 1 0 5784 0 1 -672
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1744368984
transform 1 0 3984 0 1 -672
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2
timestamp 1744368984
transform 1 0 3984 0 1 -1672
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3
timestamp 1744368984
transform 1 0 5784 0 1 -1672
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_0 JNW_ATR_SKY130A
timestamp 1744368984
transform 1 0 -1416 0 1 5528
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_1
timestamp 1744368984
transform 1 0 -1416 0 1 4128
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_2
timestamp 1744368984
transform 1 0 2184 0 1 4128
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_3
timestamp 1744368984
transform 1 0 384 0 1 6928
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_4
timestamp 1744368984
transform 1 0 3984 0 1 5528
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_5
timestamp 1744368984
transform 1 0 2184 0 1 5528
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_6
timestamp 1744368984
transform 1 0 384 0 1 5528
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_7
timestamp 1744368984
transform 1 0 384 0 1 4128
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_8
timestamp 1744368984
transform 1 0 3984 0 1 4128
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_9
timestamp 1744368984
transform 1 0 2184 0 1 6928
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_10
timestamp 1744368984
transform 1 0 3984 0 1 6928
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_11
timestamp 1744368984
transform 1 0 5784 0 1 928
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_12
timestamp 1744368984
transform 1 0 3984 0 1 928
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_13
timestamp 1744368984
transform 1 0 -1416 0 1 7028
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_14
timestamp 1744368984
transform 1 0 3984 0 1 2428
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_15
timestamp 1744368984
transform 1 0 5784 0 1 2328
box -184 -128 1336 928
use JNWTR_RPPO16  x1 JNW_TR_SKY130A
timestamp 1744468687
transform 1 0 -1000 0 1 200
box 0 0 4472 3440
use JNWTR_RPPO16  x4
timestamp 1744468687
transform -1 0 3472 0 1 -3400
box 0 0 4472 3440
use JNWATR_PCH_4C5F0  x5
timestamp 1744368984
transform 1 0 5784 0 1 5528
box -184 -128 1336 928
<< labels >>
flabel metal1 1304 8104 1496 8296 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel locali 3400 -3400 3900 -2900 0 FreeSans 1600 0 0 0 VSS
port 12 nsew
flabel metal1 6456 500 6648 692 0 FreeSans 1600 0 0 0 VOUT
port 14 nsew
flabel metal2 7136 3168 7200 3232 0 FreeSans 1600 0 0 0 VINN
port 16 nsew
flabel metal3 7134 3572 7198 3636 0 FreeSans 1600 0 0 0 VINP
port 19 nsew
<< properties >>
string FIXED_BBOX 0 0 14704 3440
<< end >>
