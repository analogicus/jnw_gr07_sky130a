magic
tech sky130A
magscale 1 2
timestamp 1744474159
<< locali >>
rect 5702 7704 9832 8100
rect 8488 7328 8680 7704
rect 9640 7376 9832 7704
rect 8488 4576 8680 6896
rect 9640 4576 9832 6996
rect 8488 3896 8680 4096
rect 9640 3896 9832 4096
rect 8488 3704 9832 3896
rect 0 3300 4500 3500
rect 4400 296 4500 3300
rect 4400 104 5396 296
rect 3868 -680 4108 20
rect 4400 0 4500 104
rect 7840 -1900 8032 -1704
rect 5000 -2000 8536 -1900
rect 4600 -2100 8536 -2000
rect 4400 -2546 8536 -2100
rect 4400 -2594 7156 -2546
rect 7204 -2594 8536 -2546
rect 4400 -2600 8536 -2594
rect 4400 -2900 9600 -2600
rect 4400 -3500 5200 -2900
rect 0 -3739 5200 -3500
rect 6100 -3739 6800 -2900
rect 7700 -3664 8400 -2900
rect 7700 -3739 8461 -3664
rect 0 -3800 5261 -3739
rect 5964 -3800 8536 -3739
rect 9300 -3800 9600 -2900
rect 0 -3900 9600 -3800
rect 0 -7100 100 -3900
rect 4400 -4500 9600 -3900
rect 4400 -5400 5261 -4500
rect 6100 -5339 6800 -4500
rect 6079 -5400 6936 -5339
rect 7700 -5400 8461 -4500
rect 9300 -5400 9600 -4500
rect 4400 -6100 9600 -5400
rect 4400 -6136 5261 -6100
rect 6064 -6121 8461 -6100
rect 4400 -7000 5200 -6136
rect 6100 -7000 6800 -6121
rect 7700 -6136 8461 -6121
rect 7700 -7000 8400 -6136
rect 9300 -7000 9600 -6100
rect 4400 -7075 9600 -7000
rect 4251 -7100 9600 -7075
rect 0 -7500 9600 -7100
rect 0 -10700 100 -7500
rect 4400 -10700 4900 -7500
rect 9200 -10700 9300 -7500
rect 0 -10800 9300 -10700
<< viali >>
rect 7156 -2594 7204 -2546
rect 364 -4280 604 -4040
rect 3880 -4280 4108 -4040
rect 380 -7880 620 -7640
rect 3868 -7880 4108 -7640
rect 5164 -7880 5404 -7640
rect 8668 -7880 8908 -7640
<< metal1 >>
rect 2274 7904 9064 8096
rect 8744 3532 8808 6932
rect 8872 4304 9064 7904
rect 9256 6404 9448 6996
rect 9256 5096 9448 5596
rect 9256 4898 9448 4904
rect 8168 3468 8808 3532
rect 9256 3696 9448 4196
rect 9256 3498 9448 3504
rect 5104 304 5476 496
rect 8168 432 8232 3468
rect 7468 368 8232 432
rect 7648 328 8232 368
rect 8168 -968 8232 328
rect 8168 -1032 8568 -968
rect 8632 -1032 8638 -968
rect 4574 -2468 4580 -2228
rect 4820 -2468 4826 -2228
rect 180 -4040 620 -4020
rect 180 -4280 364 -4040
rect 604 -4280 620 -4040
rect 180 -4300 620 -4280
rect 3874 -4040 4114 -4028
rect 4580 -4040 4820 -2468
rect 7370 -2540 7430 -2534
rect 7144 -2546 7370 -2540
rect 7144 -2594 7156 -2546
rect 7204 -2594 7370 -2546
rect 7144 -2600 7370 -2594
rect 7370 -2606 7430 -2600
rect 5800 -3180 8600 -3100
rect 5580 -3400 8908 -3180
rect 3874 -4280 3880 -4040
rect 4108 -4280 4820 -4040
rect 5400 -3600 9100 -3400
rect 3874 -4292 4114 -4280
rect 180 -7620 420 -4300
rect 5400 -6300 5900 -3600
rect 7180 -4080 7420 -4074
rect 7180 -5020 7420 -4320
rect 8600 -6300 9100 -3600
rect 5400 -6400 9100 -6300
rect 5400 -6500 8908 -6400
rect 5580 -6620 8908 -6500
rect 5900 -6800 8908 -6620
rect 8668 -7620 8908 -6800
rect 180 -7640 640 -7620
rect 180 -7880 380 -7640
rect 620 -7880 640 -7640
rect 180 -7900 640 -7880
rect 3860 -7640 4120 -7620
rect 5140 -7640 5420 -7620
rect 3860 -7880 3868 -7640
rect 4108 -7880 5164 -7640
rect 5404 -7880 5420 -7640
rect 3860 -7900 4120 -7880
rect 5140 -7900 5420 -7880
rect 8660 -7640 8920 -7620
rect 8660 -7880 8668 -7640
rect 8908 -7880 8920 -7640
rect 8660 -7900 8920 -7880
<< via1 >>
rect 9256 4904 9448 5096
rect 9256 3504 9448 3696
rect 8568 -1032 8632 -968
rect 4580 -2468 4820 -2228
rect 7370 -2600 7430 -2540
rect 7180 -4320 7420 -4080
<< metal2 >>
rect 8095 4904 8104 5096
rect 8286 4904 9256 5096
rect 9448 4904 9454 5096
rect 8080 3696 9520 3720
rect 8080 3504 9256 3696
rect 9448 3504 9520 3696
rect 8080 3480 9520 3504
rect 4580 -2228 4820 -2222
rect 4820 -2468 5950 -2228
rect 6180 -2468 6189 -2228
rect 4580 -2474 4820 -2468
rect 7632 -2540 7688 -2533
rect 7364 -2600 7370 -2540
rect 7430 -2542 7690 -2540
rect 7430 -2598 7632 -2542
rect 7688 -2598 7690 -2542
rect 7430 -2600 7690 -2598
rect 7632 -2607 7688 -2600
rect 8080 -4080 8320 3480
rect 8568 -968 8632 -962
rect 8632 -1032 8776 -968
rect 8832 -1032 8841 -968
rect 8568 -1038 8632 -1032
rect 7174 -4320 7180 -4080
rect 7420 -4320 8320 -4080
<< via2 >>
rect 8104 4904 8286 5096
rect 5950 -2468 6180 -2228
rect 7632 -2598 7688 -2542
rect 8776 -1032 8832 -968
<< metal3 >>
rect 8080 5096 8320 5120
rect 8080 4904 8104 5096
rect 8286 4904 8320 5096
rect 5945 -2228 6185 -2223
rect 8080 -2228 8320 4904
rect 8771 -968 8837 -963
rect 8768 -1032 8776 -968
rect 8832 -1032 9332 -968
rect 8771 -1037 8837 -1032
rect 9268 -1320 9332 -1032
rect 9268 -1532 9336 -1320
rect 5945 -2468 5950 -2228
rect 6180 -2468 8320 -2228
rect 5945 -2473 6185 -2468
rect 7627 -2540 7693 -2537
rect 7938 -2538 8002 -2532
rect 7627 -2542 7938 -2540
rect 7627 -2598 7632 -2542
rect 7688 -2598 7938 -2542
rect 7627 -2600 7938 -2598
rect 7627 -2603 7693 -2600
rect 7938 -2608 8002 -2602
<< via3 >>
rect 7938 -2602 8002 -2538
<< metal4 >>
rect 8400 -2400 8960 -2340
rect 7937 -2538 8003 -2537
rect 7937 -2602 7938 -2538
rect 8002 -2540 8003 -2538
rect 8400 -2540 8460 -2400
rect 8002 -2600 8460 -2540
rect 8002 -2602 8003 -2600
rect 7937 -2603 8003 -2602
use amplifier_rev2  amplifier_rev2_0 ../JNW_GR07_SKY130A
timestamp 1744468687
transform 1 0 1000 0 1 -200
box -1600 -3400 7200 8300
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1736794646
transform 1 0 8200 0 1 -5600
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1736794646
transform 1 0 5000 0 1 -7200
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1736794646
transform 1 0 5000 0 1 -5600
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1736794646
transform 1 0 6600 0 1 -7200
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1736794646
transform 1 0 8200 0 1 -7200
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1736794646
transform 1 0 5000 0 1 -4000
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1736794646
transform 1 0 6600 0 1 -4000
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1736794646
transform 1 0 6600 0 1 -5600
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1736794646
transform 1 0 8200 0 1 -4000
box 0 0 1340 1340
use JNWATR_PCH_4C5F0  x3 ../JNW_ATR_SKY130A
timestamp 1744368984
transform 1 0 8584 0 1 3928
box -184 -128 1336 928
use JNWTR_RPPO16  x4 ../JNW_TR_SKY130A
timestamp 1744468687
transform 1 0 0 0 1 -7200
box 0 0 4472 3440
use JNWATR_PCH_4C5F0  x5
timestamp 1744368984
transform 1 0 8584 0 1 6728
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  x
timestamp 1744368984
transform 1 0 8584 0 1 5328
box -184 -128 1336 928
use JNWTR_CAPX1  x2 ../JNW_TR_SKY130A
timestamp 1744368984
transform 1 0 8900 0 1 -2400
box 0 0 1080 1080
use JNWTR_RPPO16  x6
timestamp 1744468687
transform -1 0 4472 0 1 -10800
box 0 0 4472 3440
use JNWTR_RPPO16  x7
timestamp 1744468687
transform -1 0 9272 0 1 -10800
box 0 0 4472 3440
<< labels >>
flabel metal1 9256 6404 9448 6596 0 FreeSans 1600 0 0 0 I_OUT
port 1 nsew
flabel locali 4400 -10800 4900 -10300 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
flabel metal1 2304 7904 2496 8096 0 FreeSans 1600 0 0 0 VDD
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 32656 3440
<< end >>
